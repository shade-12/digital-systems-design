module tb_rtl_dotoptact();
endmodule: tb_rtl_dotoptact
