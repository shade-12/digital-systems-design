module reverse(
  input logic clk, input logic rst_n,
  input  logic [7:0] din,  input  logic din_valid,
  output logic [7:0] dout, input  logic rdy, output logic ena
);

  parameter N = 4;
  
  // your code here

endmodule
