module tb_rtl_dotopt();
endmodule: tb_rtl_dotopt
